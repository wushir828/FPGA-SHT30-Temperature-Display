module pixel_rom (
    input   wire    [8:0]   address,
    output  reg     [63:0]  q
);
    always@(*)
        case (address)
            9'd0    : q = 64'h0000000000000000;
            9'd1    : q = 64'h00000001FFE00000;
            9'd2    : q = 64'h0000001FFFFE0000;
            9'd3    : q = 64'h000000FFFFFF8000;
            9'd4    : q = 64'h000001FFFFFFE000;
            9'd5    : q = 64'h000007FFFFFFF800;
            9'd6    : q = 64'h00000FFFFFFFFC00;
            9'd7    : q = 64'h00001FF00003FE00;
            9'd8    : q = 64'h00001F0000007E00;
            9'd9    : q = 64'h00003C0000000F00;
            9'd10   : q = 64'h0000380000000700;
            9'd11   : q = 64'h0000300000000300;
            9'd12   : q = 64'h0000300000000300;
            9'd13   : q = 64'h0000300000000300;
            9'd14   : q = 64'h0000380000000700;
            9'd15   : q = 64'h0000380000000700;
            9'd16   : q = 64'h00003E0000001F00;
            9'd17   : q = 64'h00001F8000003E00;
            9'd18   : q = 64'h00001FF00003FE00;
            9'd19   : q = 64'h00000FFFFFFFFC00;
            9'd20   : q = 64'h000007FFFFFFF800;
            9'd21   : q = 64'h000003FFFFFFF000;
            9'd22   : q = 64'h000000FFFFFFC000;
            9'd23   : q = 64'h0000003FFFFF0000;
            9'd24   : q = 64'h00000003FFF00000;
            9'd25   : q = 64'h0000000000000000;
            9'd26   : q = 64'h0000000000000000;
            9'd27   : q = 64'h0000000000000000;
            9'd28   : q = 64'h0000000000000000;
            9'd29   : q = 64'h0000000000000000;
            9'd30   : q = 64'h0000000000000000;
            9'd31   : q = 64'h0000000000000000;

            9'd32   : q = 64'h0000000000000000;                
            9'd33   : q = 64'h0000000000000000;
            9'd34   : q = 64'h0000000000000000;
            9'd35   : q = 64'h0000000000000000;
            9'd36   : q = 64'h0000000000000000;
            9'd37   : q = 64'h0000000000000000;
            9'd38   : q = 64'h0000060000000300;
            9'd39   : q = 64'h0000060000000300;
            9'd40   : q = 64'h0000060000000300;
            9'd41   : q = 64'h0000060000000300;
            9'd42   : q = 64'h0000060000000300;
            9'd43   : q = 64'h0000070000000700;
            9'd44   : q = 64'h00000FFFFFFFFF00;
            9'd45   : q = 64'h00001FFFFFFFFF00;
            9'd46   : q = 64'h00003FFFFFFFFF00;
            9'd47   : q = 64'h00003FFFFFFFFF00;
            9'd48   : q = 64'h00003FFFFFFFFF00;
            9'd49   : q = 64'h0000000000000700;
            9'd50   : q = 64'h0000000000000300;
            9'd51   : q = 64'h0000000000000300;
            9'd52   : q = 64'h0000000000000300;
            9'd53   : q = 64'h0000000000000300;
            9'd54   : q = 64'h0000000000000300;
            9'd55   : q = 64'h0000000000000000;
            9'd56   : q = 64'h0000000000000000;
            9'd56   : q = 64'h0000000000000000;
            9'd57   : q = 64'h0000000000000000;
            9'd58   : q = 64'h0000000000000000;
            9'd59   : q = 64'h0000000000000000;
            9'd60   : q = 64'h0000000000000000;
            9'd61   : q = 64'h0000000000000000;
            9'd62   : q = 64'h0000000000000000;
            9'd63   : q = 64'h0000000000000000;

            9'd64   : q = 64'h00007E0000000000;
            9'd65   : q = 64'h0000000000000F00;
            9'd66   : q = 64'h000000FC00001F00;
            9'd67   : q = 64'h000003FE00007F00;
            9'd68   : q = 64'h000007FE0000FF00;
            9'd69   : q = 64'h00000FFE0001FF00;
            9'd70   : q = 64'h00001FFE0003EF00;
            9'd71   : q = 64'h00001C1E00078F00;
            9'd72   : q = 64'h00003800000F0F00;
            9'd73   : q = 64'h00003800003E0F00;
            9'd74   : q = 64'h00003000007C0F00;
            9'd75   : q = 64'h0000300000F80F00;
            9'd76   : q = 64'h0000300001F00F00;
            9'd77   : q = 64'h0000300003E00F00;
            9'd78   : q = 64'h0000300007C00F00;
            9'd79   : q = 64'h000038000F800F00;
            9'd80   : q = 64'h000038003F000F00;
            9'd81   : q = 64'h00003E00FE000F00;
            9'd82   : q = 64'h00001FC7FC000F00;
            9'd83   : q = 64'h00001FFFF8001F00;
            9'd84   : q = 64'h00000FFFF0003F00;
            9'd85   : q = 64'h000007FFC001FF00;
            9'd86   : q = 64'h000003FF8003FF00;
            9'd87   : q = 64'h0000007C0003F000;
            9'd88   : q = 64'h0000000000000000;
            9'd89   : q = 64'h0000000000000000;
            9'd90   : q = 64'h0000000000000000;
            9'd91   : q = 64'h0000000000000000;
            9'd92   : q = 64'h0000000000000000;
            9'd93   : q = 64'h0000000000000000;
            9'd94   : q = 64'h0000000000000000;
            9'd95   : q = 64'h0000000000000000;

            9'd96   : q = 64'h0000000000000000;
            9'd97   : q = 64'h0000000000000000; 
            9'd98   : q = 64'h000000E00003F000; 
            9'd99   : q = 64'h000003F00003F800; 
            9'd100  : q = 64'h00000FF80007FC00; 
            9'd101  : q = 64'h00000FF80007FE00; 
            9'd102  : q = 64'h00001FF80003FE00; 
            9'd103  : q = 64'h00001C700003CF00; 
            9'd104  : q = 64'h0000380000000700; 
            9'd105  : q = 64'h0000300018000300; 
            9'd106  : q = 64'h0000300018000300; 
            9'd107  : q = 64'h0000300038000300; 
            9'd108  : q = 64'h0000300038000300; 
            9'd109  : q = 64'h0000300038000300; 
            9'd110  : q = 64'h000038007C000300; 
            9'd111  : q = 64'h000038007C000700; 
            9'd112  : q = 64'h00003E00FE000F00; 
            9'd113  : q = 64'h00001FFFEF001E00; 
            9'd114  : q = 64'h00001FFFEFC07E00; 
            9'd115  : q = 64'h00000FFFC7FFFC00; 
            9'd116  : q = 64'h000007FF83FFFC00;  
            9'd117  : q = 64'h000003FE01FFF800; 
            9'd118  : q = 64'h0000007800FFE000; 
            9'd119  : q = 64'h00000000003F8000; 
            9'd120  : q = 64'h0000000000000000; 
            9'd121  : q = 64'h0000000000000000; 
            9'd122  : q = 64'h0000000000000000; 
            9'd123  : q = 64'h0000000000000000; 
            9'd124  : q = 64'h0000000000000000; 
            9'd125  : q = 64'h0000000000000000; 
            9'd126  : q = 64'h0000000000000000; 
            9'd127  : q = 64'h0000000000000000; 

            9'd128  : q = 64'h0000000000000000;
            9'd129  : q = 64'h0000000000180000;
            9'd130  : q = 64'h0000000000780000;
            9'd131  : q = 64'h0000000001F80000;
            9'd132  : q = 64'h0000000003F80000;
            9'd133  : q = 64'h000000000FD80000;
            9'd134  : q = 64'h000000001F180000;
            9'd135  : q = 64'h000000007E180000;
            9'd136  : q = 64'h00000000F8180000;
            9'd137  : q = 64'h00000003E0180000;
            9'd138  : q = 64'h0000000FC0180300;
            9'd139  : q = 64'h0000001F00180300;
            9'd140  : q = 64'h0000007E00180300;
            9'd141  : q = 64'h000000F800180300;
            9'd142  : q = 64'h000003E000180300;
            9'd143  : q = 64'h000007C000180700;
            9'd144  : q = 64'h00001FFFFFFFFF00;
            9'd145  : q = 64'h00003FFFFFFFFF00;
            9'd146  : q = 64'h00003FFFFFFFFF00;
            9'd147  : q = 64'h00003FFFFFFFFF00;
            9'd148  : q = 64'h00003FFFFFFFFF00;
            9'd149  : q = 64'h0000000000180300;
            9'd150  : q = 64'h0000000000180300;
            9'd151  : q = 64'h0000000000180300;
            9'd152  : q = 64'h0000000000180300;
            9'd153  : q = 64'h0000000000180300;
            9'd154  : q = 64'h0000000000180000;
            9'd155  : q = 64'h0000000000000000;
            9'd156  : q = 64'h0000000000000000;
            9'd157  : q = 64'h0000000000000000;
            9'd158  : q = 64'h0000000000000000;
            9'd159  : q = 64'h0000000000000000;

            9'd160  : q = 64'h0000000000000000;
            9'd161  : q = 64'h0000000000000000;
            9'd162  : q = 64'h000000000003E000;
            9'd163  : q = 64'h00000001FC07F800;
            9'd164  : q = 64'h00003FFFFC0FFC00;
            9'd165  : q = 64'h00003FFFFC0FFC00;
            9'd166  : q = 64'h00003FFFFC07FE00;
            9'd167  : q = 64'h00003C0078078600;
            9'd168  : q = 64'h00003C00F0000700;
            9'd169  : q = 64'h00003C00E0000300;
            9'd170  : q = 64'h00003C01C0000300;
            9'd171  : q = 64'h00003C01C0000300;
            9'd172  : q = 64'h00003C01C0000300;
            9'd173  : q = 64'h00003C01C0000300;
            9'd174  : q = 64'h00003C01C0000300;
            9'd175  : q = 64'h00003C01E0000700;
            9'd176  : q = 64'h00003C01E0000F00;
            9'd177  : q = 64'h00003C00F8001F00;
            9'd178  : q = 64'h00003C00FE00FE00;
            9'd179  : q = 64'h00003C00FFFFFE00;
            9'd180  : q = 64'h00003C007FFFFC00;
            9'd181  : q = 64'h00003C003FFFF800;
            9'd182  : q = 64'h000038000FFFE000;
            9'd183  : q = 64'h0000200003FF8000;
            9'd184  : q = 64'h0000000000000000;
            9'd185  : q = 64'h0000000000000000;
            9'd186  : q = 64'h0000000000000000;
            9'd187  : q = 64'h0000000000000000;
            9'd188  : q = 64'h0000000000000000;
            9'd189  : q = 64'h0000000000000000;
            9'd190  : q = 64'h0000000000000000;
            9'd191  : q = 64'h0000000000000000;

            9'd192  : q = 64'h0000000000000000;
            9'd193  : q = 64'h0000000000000000;
            9'd194  : q = 64'h0000000000000000;
            9'd195  : q = 64'h0000000000000000;
            9'd196  : q = 64'h00000001FFF80000;
            9'd197  : q = 64'h0000001FFFFF8000;
            9'd198  : q = 64'h0000007FFFFFE000;
            9'd199  : q = 64'h000001FFFFFFF000;
            9'd200  : q = 64'h000003FFFFFFF800;
            9'd201  : q = 64'h000007FFFFFFFC00;
            9'd202  : q = 64'h00000FE03E00FE00;
            9'd203  : q = 64'h00001F0078003E00;
            9'd204  : q = 64'h00001E0070000F00;
            9'd205  : q = 64'h00003C00F0000700;
            9'd206  : q = 64'h00003800E0000700;
            9'd207  : q = 64'h00003000E0000300;
            9'd208  : q = 64'h00003001C0000300;
            9'd209  : q = 64'h00003001C0000300;
            9'd210  : q = 64'h00003001E0000300;
            9'd211  : q = 64'h00003000E0000700;
            9'd212  : q = 64'h00003F80F0000F00;
            9'd213  : q = 64'h00003FC0FC001E00;
            9'd214  : q = 64'h00003FC0FF83FE00;
            9'd215  : q = 64'h00001FC07FFFFC00;
            9'd216  : q = 64'h00000F803FFFF800;
            9'd217  : q = 64'h000007801FFFF000;
            9'd218  : q = 64'h0000000007FFC000;
            9'd219  : q = 64'h0000000000FE0000;
            9'd220  : q = 64'h0000000000000000;
            9'd221  : q = 64'h0000000000000000;
            9'd222  : q = 64'h0000000000000000;
            9'd223  : q = 64'h0000000000000000;

            9'd224  : q = 64'h0000000000000000;
            9'd225  : q = 64'h0000000000000000;
            9'd226  : q = 64'h0000000000000000;
            9'd227  : q = 64'h0000000000000000;
            9'd228  : q = 64'h000001F000000000;
            9'd229  : q = 64'h00003FF000000000;
            9'd230  : q = 64'h00003FE000000000;
            9'd231  : q = 64'h00003F0000000000;
            9'd232  : q = 64'h00003E0000000000;
            9'd233  : q = 64'h00003C0000000000;
            9'd234  : q = 64'h00003C000000FE00;
            9'd235  : q = 64'h00003C00000FFF00;
            9'd236  : q = 64'h00003C0000FFFF00;
            9'd237  : q = 64'h00003C0003FFFF00;
            9'd238  : q = 64'h00003C000FFFFF00;
            9'd239  : q = 64'h00003C007FFFFF00;
            9'd240  : q = 64'h00003C01FFF8FC00;
            9'd241  : q = 64'h00003C07FE000000;
            9'd242  : q = 64'h00003C1FF0000000;
            9'd243  : q = 64'h00003C3F80000000;
            9'd244  : q = 64'h00003CFE00000000;
            9'd245  : q = 64'h00003FF800000000;
            9'd246  : q = 64'h00003FE000000000;
            9'd247  : q = 64'h00003F8000000000;
            9'd248  : q = 64'h00003E0000000000;
            9'd249  : q = 64'h0000380000000000;
            9'd250  : q = 64'h0000000000000000;
            9'd251  : q = 64'h0000000000000000;
            9'd252  : q = 64'h0000000000000000;
            9'd253  : q = 64'h0000000000000000;
            9'd254  : q = 64'h0000000000000000;
            9'd255  : q = 64'h0000000000000000;

            9'd256  : q = 64'h0000000000000000;
            9'd257  : q = 64'h0000000000000000;
            9'd258  : q = 64'h0000000000000000;
            9'd259  : q = 64'h0000000000000000;
            9'd260  : q = 64'h000000FC003FC000;
            9'd261  : q = 64'h000003FF00FFF000;
            9'd262  : q = 64'h000007FF81FFF800;
            9'd263  : q = 64'h00000FFFC3FFFC00;
            9'd264  : q = 64'h00001FFFE7FCFE00;
            9'd265  : q = 64'h00001E01EFE01E00;
            9'd266  : q = 64'h00003C00FFC00F00;
            9'd267  : q = 64'h000038007F800700;
            9'd268  : q = 64'h000030003F000300;
            9'd269  : q = 64'h000030003F000300;
            9'd270  : q = 64'h000030003E000300;
            9'd271  : q = 64'h000030007C000300;
            9'd272  : q = 64'h000030007C000300;
            9'd273  : q = 64'h00003000F8000300;
            9'd274  : q = 64'h00003800FC000700;
            9'd275  : q = 64'h00003801FE000700;
            9'd276  : q = 64'h00001C03FF000E00;
            9'd277  : q = 64'h00001F0FEF801E00;
            9'd278  : q = 64'h00000FFFC7F07C00;
            9'd279  : q = 64'h00000FFFC3FFFC00;
            9'd280  : q = 64'h000003FF01FFF800;
            9'd281  : q = 64'h000001FE00FFF000;
            9'd282  : q = 64'h00000000003FC000;
            9'd283  : q = 64'h0000000000000000;
            9'd284  : q = 64'h0000000000000000;
            9'd285  : q = 64'h0000000000000000;
            9'd286  : q = 64'h0000000000000000;
            9'd287  : q = 64'h0000000000000000;

            9'd288  : q = 64'h0000000000000000;
            9'd289  : q = 64'h0000000000000000;
            9'd290  : q = 64'h0000007FF0000000;
            9'd291  : q = 64'h000001FFFC000000;
            9'd292  : q = 64'h000003FFFE007C00;
            9'd293  : q = 64'h00000FFFFF00FE00;
            9'd294  : q = 64'h00000FFFFF80FE00;
            9'd295  : q = 64'h00001F803F80FF00;
            9'd296  : q = 64'h00003E0007C07F00;
            9'd297  : q = 64'h0000380003C03F00;
            9'd298  : q = 64'h0000380001C00300;
            9'd299  : q = 64'h0000300001C00300;
            9'd300  : q = 64'h0000300001C00300;
            9'd301  : q = 64'h0000300001C00300;
            9'd302  : q = 64'h0000300001C00700;
            9'd303  : q = 64'h0000300003C00F00;
            9'd304  : q = 64'h0000380003801E00;
            9'd305  : q = 64'h00003C0007807E00;
            9'd306  : q = 64'h00001E001F01FC00;
            9'd307  : q = 64'h00001FC07E3FF800;
            9'd308  : q = 64'h00000FFFFFFFF000;
            9'd309  : q = 64'h000007FFFFFFE000;
            9'd310  : q = 64'h000003FFFFFF8000;
            9'd311  : q = 64'h000000FFFFFE0000;
            9'd312  : q = 64'h0000003FFFF00000;
            9'd313  : q = 64'h00000001FE000000;
            9'd314  : q = 64'h0000000000000000;
            9'd315  : q = 64'h0000000000000000;
            9'd316  : q = 64'h0000000000000000;
            9'd317  : q = 64'h0000000000000000;
            9'd318  : q = 64'h0000000000000000;
            9'd319  : q = 64'h0000000000000000;

            9'd320  : q = 64'h0000000000000000;
            9'd321  : q = 64'h000FFFFFFFFFFF80;
            9'd322  : q = 64'h000FFFFFFFFFFF80;
            9'd323  : q = 64'h000FFFFFFFFFFF80;
            9'd324  : q = 64'h000FFFFFFFFFFF80;
            9'd325  : q = 64'h000FFFFFFFFFFF80;
            9'd326  : q = 64'h000FFFFFFFFFFF80;
            9'd327  : q = 64'h00000000F8000000;
            9'd328  : q = 64'h00000000F8000000;
            9'd329  : q = 64'h00000000F8000000;
            9'd330  : q = 64'h00000000F8000000;
            9'd331  : q = 64'h00000000F8000000;
            9'd332  : q = 64'h00000000F8000000;
            9'd333  : q = 64'h00000000F8000000;
            9'd334  : q = 64'h00000000F8000000;
            9'd335  : q = 64'h00000000F8000000;
            9'd336  : q = 64'h00000000F8000000;
            9'd337  : q = 64'h00000000F8000000;
            9'd338  : q = 64'h00000000F8000000;
            9'd339  : q = 64'h00000000F8000000;
            9'd340  : q = 64'h00000000F8000000;
            9'd341  : q = 64'h00000000F8000000;
            9'd342  : q = 64'h00000000F8000000;
            9'd343  : q = 64'h00000000F8000000;
            9'd344  : q = 64'h000FFFFFFFFFFF80;
            9'd345  : q = 64'h000FFFFFFFFFFF80;
            9'd346  : q = 64'h000FFFFFFFFFFF80;
            9'd347  : q = 64'h000FFFFFFFFFFF80;
            9'd348  : q = 64'h000FFFFFFFFFFF80;
            9'd349  : q = 64'h000FFFFFFFFFFF80;
            9'd350  : q = 64'h0000000000000000;
            9'd351  : q = 64'h0000000000000000;

            9'd352  : q = 64'h0000000000000000;
            9'd353  : q = 64'h0007E00000000000;
            9'd354  : q = 64'h0007E00000000000;
            9'd355  : q = 64'h0007E00000000000;
            9'd356  : q = 64'h0007E00000000000;
            9'd357  : q = 64'h0007E00000000000;
            9'd358  : q = 64'h0007E00000000000;
            9'd359  : q = 64'h0007E00000000000;
            9'd360  : q = 64'h0007E00000000000;
            9'd361  : q = 64'h0007E00000000000;
            9'd362  : q = 64'h0007E00000000000;
            9'd363  : q = 64'h0007E00000000000;
            9'd364  : q = 64'h0007FFFFFFFFFF00;
            9'd365  : q = 64'h0007FFFFFFFFFF00;
            9'd366  : q = 64'h0007FFFFFFFFFF00;
            9'd367  : q = 64'h0007FFFFFFFFFF00;
            9'd368  : q = 64'h0007FFFFFFFFFF00;
            9'd369  : q = 64'h0007FFFFFFFFFF00;
            9'd370  : q = 64'h0007FFFFFFFFFF00;
            9'd371  : q = 64'h0007E00000000000;
            9'd372  : q = 64'h0007E00000000000;
            9'd373  : q = 64'h0007E00000000000;
            9'd374  : q = 64'h0007E00000000000;
            9'd375  : q = 64'h0007E00000000000;
            9'd376  : q = 64'h0007E00000000000;
            9'd377  : q = 64'h0007E00000000000;
            9'd378  : q = 64'h0007E00000000000;
            9'd379  : q = 64'h0007E00000000000;
            9'd380  : q = 64'h0007E00000000000;
            9'd381  : q = 64'h0007E00000000000;
            9'd382  : q = 64'h0007E00000000000;
            9'd383  : q = 64'h0003E00000000000;
            9'd384  : q = 64'h0000000000000000;
            //-
            9'd385  : q = 64'h0000000000000000;
            9'd386  : q = 64'h0000000000000000;
            9'd387  : q = 64'h0000000000000000;
            9'd388  : q = 64'h0000000000000000;
            9'd389  : q = 64'h0000000000000000;
            9'd390  : q = 64'h000000003c000000;
            9'd391  : q = 64'h000000003c000000;
            9'd392  : q = 64'h000000003c000000;
            9'd393  : q = 64'h000000003c000000;
            9'd394  : q = 64'h000000003c000000;
            9'd395  : q = 64'h000000003c000000;
            9'd396  : q = 64'h000000003c000000;
            9'd397  : q = 64'h000000003c000000;
            9'd398  : q = 64'h000000003c000000; 
            9'd399  : q = 64'h000000003c000000; 
            9'd400  : q = 64'h000000003c000000; 
            9'd401  : q = 64'h000000003c000000; 
            9'd402  : q = 64'h000000003c000000; 
            9'd403  : q = 64'h000000003c000000; 
            9'd404  : q = 64'h000000003c000000; 
            9'd405  : q = 64'h000000003c000000; 
            9'd406  : q = 64'h000000003c000000; 
            9'd407  : q = 64'h000000003c000000; 
            9'd408  : q = 64'h000000003c000000; 
            9'd409  : q = 64'h000000003c000000; 
            9'd410  : q = 64'h0000000000000000;
            9'd411  : q = 64'h0000000000000000;
            9'd412  : q = 64'h0000000000000000;
            9'd413  : q = 64'h0000000000000000;
            9'd414  : q = 64'h0000000000000000;
            9'd415  : q = 64'h0000000000000000;
            9'd416  : q = 64'h0000000000000000;
            9'd417  : q = 64'h0000000000000000;
            //.
            9'd418  : q = 64'h0000000000000000;
            9'd419  : q = 64'h000000000000ff00;
            9'd420  : q = 64'h000000000000ff00;
            9'd421  : q = 64'h000000000000ff00;
            9'd422  : q = 64'h000000000000ff00;
            9'd423  : q = 64'h000000000000ff00;
            9'd424  : q = 64'h000000000000ff00;
            9'd425  : q = 64'h000000000000ff00;
            9'd426  : q = 64'h000000000000ff00;
            9'd427  : q = 64'h0000000000000000;
            9'd428  : q = 64'h0000000000000000;
            9'd429  : q = 64'h0000000000000000;
        //:
            9'd430  : q = 64'h0000000000000000;
            9'd431  : q = 64'h0000000001801C00;
            9'd432  : q = 64'h0000000007E03F00;
            9'd433  : q = 64'h000000000FF07F80;
            9'd434  : q = 64'h000000000FF07F80;
            9'd435  : q = 64'h000000000FF07F80;
            9'd436  : q = 64'h000000000FF07F80;
            9'd437  : q = 64'h000000000FF07F80;
            9'd438  : q = 64'h000000000FF07F80;
            9'd439  : q = 64'h0000000007E03F00;
            9'd440  : q = 64'h0000000003C00C00;
            9'd441  : q = 64'h0000000000000000;
            9'd442  : q = 64'h0000000000000000;
            default: q = 16'h0;
        endcase
endmodule